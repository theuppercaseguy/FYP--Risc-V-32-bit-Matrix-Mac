module gate(A,B,Y);
    //declare inputs
    input A,B;
    output Y;

    //gatelevel modeling
    //example
    //functionname (port list)
    //              (outputs,inputs)
    and (Y,A,B);
    


endmodule